module tb3

reg   [

